module displays;
    initial 
        begin
            $display("test");
        end
endmodule