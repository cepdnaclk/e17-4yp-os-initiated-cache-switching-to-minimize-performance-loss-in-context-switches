`include "../modules/32bit-Int-Mul/mul.v"
module testmul;


  reg [31:0] data1,data2;
  reg [2:0] select;
  wire [31:0] result;

  //cpu module instantiate RESULT, DATA1, DATA2, SELECT
  mul mymul(result, data1, data2, select);

	//wavedata file
	initial
	begin
		$dumpfile("wavedata.vcd");
		$dumpvars(0,testmul);
			
	end

	//running
	initial
	begin

		data1 = 32'b00000000000000000000000000000011;
    data2 = 32'b00000000000000000000000000000001;
    select = 3'b000;
		#1

    data1 = 32'b00000000000000000000000000000011;
    data2 = 32'b00000000000000000000000000000001;
    select = 3'b001;
		#1
    data1 = 32'b00000000000000000000000000000011;
    data2 = 32'b00000000000000000000000000000001;
    select = 3'b010;
		#1
    data1 = 32'b00000000000000000000000000000011;
    data2 = 32'b00000000000000000000000000000001;
    select = 3'b011;
		#1
    data1 = 32'b00000000000000000000000000000011;
    data2 = 32'b00000000000000000000000000000001;
    select = 3'b100;
		#1
    data1 = 32'b00000000000000000000000000000011;
    data2 = 32'b00000000000000000000000000000001;
    select = 3'b101;
		#1
    data1 = 32'b00000000000000000000000000000011;
    data2 = 32'b00000000000000000000000000000001;
    select = 3'b110;
		#1
    data1 = 32'b00000000000000000000000000000011;
    data2 = 32'b00000000000000000000000000000001;
    select = 3'b111;
		#1

    //- values

    data1 = 32'b00000000000000000000000000000011;
    data2 = 32'b11111111111111111111111111111111;
    select = 3'b000;
		#1

    data1 = 32'b00000000000000000000000000000001;
    data2 = 32'b11111111111111111111111111111111;
    select = 3'b001;
		#1

    data1 = 32'b00000000000000000000000000000001;
    data2 = 32'b11111111111111111111111111111111;
    select = 3'b010;
		#1

    data1 = 32'b11111111111111111111111111111111;
    data2 = 32'b00000000000000000000000000000001;
    select = 3'b011;
		#1

    data1 = 32'b00000000000000000000000000000011;
    data2 = 32'b11111111111111111111111111111110;
    select = 3'b011;
		#1

		$finish;

	end
			 
endmodule