module Data_load_controller (
    func3,
    data_mem_in,
    data_out
);

input [2:0] func3;
input [31:0] data_mem_in;
output reg [31:0] data_out;
wire [31:0] lb,lbu,lh,lhu;

/*
| imm[11:0] |   rs1   | 000 |  rd | 0000011 |   LB  
| imm[11:0] |   rs1   | 001 |  rd | 0000011 |   LH  
| imm[11:0] |   rs1   | 010 |  rd | 0000011 |   LW  
| imm[11:0] |   rs1   | 100 |  rd | 0000011 |   LBU 
| imm[11:0] |   rs1   | 101 |  rd | 0000011 |   LHU 
*/

assign lb ={{24{data_mem_in[7]}},data_mem_in[7:0]};
assign lbu ={{24{1'b0}},data_mem_in[7:0]};
assign lh ={{16{data_mem_in[15]}},data_mem_in[15:0]};
assign lhu ={{16{1'b0}},data_mem_in[15:0]};


always @(*) begin
    case(func3)
        3'b000:begin
            data_out<=lb;
        end
        3'b001:begin
            data_out<=lh;
        end
        3'b010:begin
            data_out<=data_mem_in;
        end
        3'b100:begin
            data_out<=lbu;
        end
        default:begin
            data_out<=lhu;
        end
    endcase
end
    
endmodule